module bf_class (
    input [15:0] a,
    output zero,
    output infinity,
    output nan,
    output
);
    
endmodule